
module UART(





);
endmodule;
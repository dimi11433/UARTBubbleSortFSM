`include uart_Receiver.v
`include uart_Transmitter.v



module UART(
    input i_CLOCK,
    input i_Rx_Serial,
    output i_Tx_Serial
);
    
    

    

endmodule;
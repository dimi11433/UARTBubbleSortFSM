
module UART(





);


endmodule;